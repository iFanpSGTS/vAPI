module attack

import discord
import os

pub fn send_attack(username string, host string, port string, times string, method string) {
	"not done yet"
	//discord.send_attack_logs(username, host, port, times, method)
}